//Subject:     CO project 2 - Adder
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:     110550148
//----------------------------------------------
//Date: 	  05/01        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Adder(
    src1_i,
	src2_i,
	sum_o
	);
     
//I/O ports
input  [32-1:0]  src1_i;
input  [32-1:0]	 src2_i;
output [32-1:0]	 sum_o;

//Internal Signals
//wire    [32-1:0]	 sum_o;
wire zero_o;
//Parameter
    
//Main function
ALU adder1(src1_i, src2_i, 4'b0010, sum_o, zero_o);
endmodule





                    
                    